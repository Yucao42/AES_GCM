
    aes_signal_passing pass0
    (
        .clk(clk),
        .i_plain_text(bytext0),
        .i_aad(byaad0),
        .i_signal(bysig0),
        .i_instance_size(byins0),
        .o_instance_size(byins1),
        .o_aad(byaad1),
        .o_signal(bysig1),
        .o_plain_text(bypass1)
    )
        
    aes_signal_passing pass1
    (
        .clk(clk),
        .i_plain_text(bytext1),
        .i_aad(byaad1),
        .i_signal(bysig1),
        .i_instance_size(byins1),
        .o_instance_size(byins2),
        .o_aad(byaad2),
        .o_signal(bysig2),
        .o_plain_text(bypass2)
    )
        
    aes_signal_passing pass2
    (
        .clk(clk),
        .i_plain_text(bytext2),
        .i_aad(byaad2),
        .i_signal(bysig2),
        .i_instance_size(byins2),
        .o_instance_size(byins3),
        .o_aad(byaad3),
        .o_signal(bysig3),
        .o_plain_text(bypass3)
    )
        
    aes_signal_passing pass3
    (
        .clk(clk),
        .i_plain_text(bytext3),
        .i_aad(byaad3),
        .i_signal(bysig3),
        .i_instance_size(byins3),
        .o_instance_size(byins4),
        .o_aad(byaad4),
        .o_signal(bysig4),
        .o_plain_text(bypass4)
    )
        
    aes_signal_passing pass4
    (
        .clk(clk),
        .i_plain_text(bytext4),
        .i_aad(byaad4),
        .i_signal(bysig4),
        .i_instance_size(byins4),
        .o_instance_size(byins5),
        .o_aad(byaad5),
        .o_signal(bysig5),
        .o_plain_text(bypass5)
    )
        
    aes_signal_passing pass5
    (
        .clk(clk),
        .i_plain_text(bytext5),
        .i_aad(byaad5),
        .i_signal(bysig5),
        .i_instance_size(byins5),
        .o_instance_size(byins6),
        .o_aad(byaad6),
        .o_signal(bysig6),
        .o_plain_text(bypass6)
    )
        
    aes_signal_passing pass6
    (
        .clk(clk),
        .i_plain_text(bytext6),
        .i_aad(byaad6),
        .i_signal(bysig6),
        .i_instance_size(byins6),
        .o_instance_size(byins7),
        .o_aad(byaad7),
        .o_signal(bysig7),
        .o_plain_text(bypass7)
    )
        
    aes_signal_passing pass7
    (
        .clk(clk),
        .i_plain_text(bytext7),
        .i_aad(byaad7),
        .i_signal(bysig7),
        .i_instance_size(byins7),
        .o_instance_size(byins8),
        .o_aad(byaad8),
        .o_signal(bysig8),
        .o_plain_text(bypass8)
    )
        
    aes_signal_passing pass8
    (
        .clk(clk),
        .i_plain_text(bytext8),
        .i_aad(byaad8),
        .i_signal(bysig8),
        .i_instance_size(byins8),
        .o_instance_size(byins9),
        .o_aad(byaad9),
        .o_signal(bysig9),
        .o_plain_text(bypass9)
    )
        
    aes_signal_passing pass9
    (
        .clk(clk),
        .i_plain_text(bytext9),
        .i_aad(byaad9),
        .i_signal(bysig9),
        .i_instance_size(byins9),
        .o_instance_size(byins10),
        .o_aad(byaad10),
        .o_signal(bysig10),
        .o_plain_text(bypass10)
    )
        
    aes_signal_passing pass10
    (
        .clk(clk),
        .i_plain_text(bytext10),
        .i_aad(byaad10),
        .i_signal(bysig10),
        .i_instance_size(byins10),
        .o_instance_size(byins11),
        .o_aad(byaad11),
        .o_signal(bysig11),
        .o_plain_text(bypass11)
    )
        
    aes_signal_passing pass11
    (
        .clk(clk),
        .i_plain_text(bytext11),
        .i_aad(byaad11),
        .i_signal(bysig11),
        .i_instance_size(byins11),
        .o_instance_size(byins12),
        .o_aad(byaad12),
        .o_signal(bysig12),
        .o_plain_text(bypass12)
    )
        
    aes_signal_passing pass12
    (
        .clk(clk),
        .i_plain_text(bytext12),
        .i_aad(byaad12),
        .i_signal(bysig12),
        .i_instance_size(byins12),
        .o_instance_size(byins13),
        .o_aad(byaad13),
        .o_signal(bysig13),
        .o_plain_text(bypass13)
    )
        
    aes_signal_passing pass13
    (
        .clk(clk),
        .i_plain_text(bytext13),
        .i_aad(byaad13),
        .i_signal(bysig13),
        .i_instance_size(byins13),
        .o_instance_size(byins14),
        .o_aad(byaad14),
        .o_signal(bysig14),
        .o_plain_text(bypass14)
    )
        
    aes_signal_passing pass14
    (
        .clk(clk),
        .i_plain_text(bytext14),
        .i_aad(byaad14),
        .i_signal(bysig14),
        .i_instance_size(byins14),
        .o_instance_size(byins15),
        .o_aad(byaad15),
        .o_signal(bysig15),
        .o_plain_text(bypass15)
    )
        